//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Mon Mar 31 15:22:45 2025
// Version: 2024.1 2024.1.0.3
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// exemploISP
module exemploISP(
    // Outputs
    o_LED
);

//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output [1:0] o_LED;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   [1:0] o_LED_net_0;
wire         OSC_C1_0_RCOSC_1MHZ_O2F;
wire   [1:0] o_LED_net_1;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire         VCC_net;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign VCC_net = 1'b1;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign o_LED_net_1 = o_LED_net_0;
assign o_LED[1:0]  = o_LED_net_1;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------led_blink
led_blink led_blink_0(
        // Inputs
        .clk    ( OSC_C1_0_RCOSC_1MHZ_O2F ),
        .resetN ( VCC_net ),
        // Outputs
        .o_LED  ( o_LED_net_0 ) 
        );

//--------OSC_C1
OSC_C1 OSC_C1_0(
        // Outputs
        .RCOSC_1MHZ_O2F ( OSC_C1_0_RCOSC_1MHZ_O2F ) 
        );


endmodule
